/*!
 * @author radigast
 */

package lab_test_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"
    
    import dstream_pkg::*;
    import a_layer_pkg::*;
    import cam_ral_pkg::*;

    `include "lab_env_config.svh"
    `include "lab_env.svh"
    `include "lab_test_example.svh"

endpackage
