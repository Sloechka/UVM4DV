/**
 * @author radigast
 */

`ifndef CAM_RAL_PKG__SV
`define CAM_RAL_PKG__SV

package cam_ral_pkg;

  `include "uvm_macros.svh"
  import uvm_pkg::*;

  `include "cam_regs.svh"
  `include "cam_reg_env.svh"

endpackage: cam_ral_pkg

`endif // CAM_RAL_PKG__SV

