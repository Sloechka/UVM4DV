typedef uvm_sequencer#(axis_transaction) axis_sequencer;
