package axis_agent_pkg;
        
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "axis_config.svh"
    `include "axis_transaction.svh"
    `include "axis_sequencer.svh"
    `include "axis_driver.svh"
    `include "axis_monitor.svh"
    `include "axis_agent.svh"

endpackage: axis_agent_pkg
