package reset_agent_pkg;
        
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "reset_config.svh"
    `include "reset_driver.svh"
    `include "reset_agent.svh"

endpackage: reset_agent_pkg
