/*!
 * @author radigast
 */

package test_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"
        
    `include "my_comps_and_objs.svh"
    `include "env.svh"
    `include "test_example.svh"

endpackage
