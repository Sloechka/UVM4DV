`timescale 1ps/1ps

interface reset_if();

    logic rst_n;

endinterface: reset_if
