package test_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"
        
    import reset_agent_pkg::*;
    import axis_agent_pkg::*;

    `include "axis_sequence.svh"
    `include "env.svh"
    `include "test.svh"

endpackage: test_pkg
